`ifndef R0
  `define R0 3'b000
`endif

`ifndef R1
  `define R1 3'b001
`endif

`ifndef R2
  `define R2 3'b010
`endif

`ifndef R3
  `define R3 3'b011
`endif

`ifndef R4
  `define R4 3'b100
`endif

`ifndef R5
  `define R5 3'b101
`endif

`ifndef R6
  `define R6 3'b110
`endif

`ifndef R7
  `define R7 3'b111
`endif
